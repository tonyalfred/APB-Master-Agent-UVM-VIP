/**********************************************************************************************************************
 *  FILE DESCRIPTION
 *  -------------------------------------------------------------------------------------------------------------------
 *  File:         apb_driver.sv
 *
 *  Description:  
 * 
 *********************************************************************************************************************/

  `ifndef APB_DRIVER
    `define APB_DRIVER

    class apb_driver extends uvm_driver #(apb_seq_item);
      `uvm_component_utils(apb_driver)

      apb_seq_item m_item;

      apb_agent_config m_cfg;
      virtual apb_if m_vif;

      function new(string name = "apb_driver", uvm_component parent = null);
        super.new(name,parent);
      endfunction

      function void build_phase (uvm_phase phase);
        super.build_phase(phase);

        if(!(uvm_config_db#(apb_agent_config)::get(this,"","apb_agent_cfg",m_cfg)))
          `uvm_fatal(get_full_name(),"Error! apb_driver failed to receive m_cfg.")
        
        `uvm_info("BUILD_PHASE", "apb_driver.", UVM_HIGH)
      endfunction

      function void connect_phase (uvm_phase phase);
        super.connect_phase(phase);

        m_vif = m_cfg.m_vif;

        `uvm_info("CONNECT_PHASE", "apb_driver.", UVM_HIGH)
      endfunction

      task run_phase (uvm_phase phase);
        super.run_phase(phase);
        `uvm_info("RUN_PHASE", "apb_driver.", UVM_HIGH)
        
        forever begin
          seq_item_port.get_next_item(m_item);
          drive_transaction(m_item);
          seq_item_port.item_done();
        end
      endtask

      task drive_transaction(apb_seq_item item);
        m_vif.cb.PADDR   <= item.m_addr;
        m_vif.cb.PWRITE  <= bit'(item.m_txn);
        m_vif.cb.PSEL    <= 1'b1;
        m_vif.cb.PENABLE <= 1'b0;

        if (item.m_txn == WRITE) begin
          m_vif.cb.PWDATA <= item.m_data;
        end

        @ (m_vif.cb)
        m_vif.cb.PENABLE <= 1'b1;

        @ (m_vif.cb)
        wait (m_vif.cb.PREADY);
        m_vif.cb.PENABLE <= 1'b0;
        m_vif.cb.PSEL    <= 1'b0;
      endtask
    endclass 
  `endif

/**********************************************************************************************************************
*  END OF FILE: apb_driver.sv
*********************************************************************************************************************/