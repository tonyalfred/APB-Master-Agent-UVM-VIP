/**********************************************************************************************************************
 *  FILE DESCRIPTION
 *  -------------------------------------------------------------------------------------------------------------------
 *  File:         apb_types.sv
 *
 *  Description:  
 * 
 *********************************************************************************************************************/

  `ifndef APB_TYPES
    `define APB_TYPES

    typedef virtual apb_if apb_vif_t;
      
    typedef enum {READ = 0, WRITE = 1} apb_transaction_type_t;

    typedef logic [`APB_DATA_WIDTH-1:0] apb_data_t;

    typedef logic [`APB_ADDR_WIDTH-1:0] apb_addr_t;
  `endif

/**********************************************************************************************************************
*  END OF FILE: apb_types.sv
*********************************************************************************************************************/