/**********************************************************************************************************************
 *  FILE DESCRIPTION
 *  -------------------------------------------------------------------------------------------------------------------
 *  File:         apb_pkg.sv
 *
 *  Description:  
 * 
 *********************************************************************************************************************/

    `include "apb_defines.sv"
    `include "apb_if.sv"

    package apb_pkg;
        import uvm_pkg::*;
        `include "uvm_macros.svh"

        `include "apb_types.sv"
        `include "apb_seq_item.sv"
        `include "apb_reset_item.sv"
        `include "apb_seq_lib.sv"
        `include "apb_virtual_seq.sv"

        `include "apb_agent_config.sv"
        `include "apb_sequencer.sv"
        `include "apb_driver.sv"
        `include "apb_monitor.sv"
        `include "apb_subscriber.sv"
        `include "apb_agent.sv"

        `include "apb_reset_sequencer.sv"
        `include "apb_reset_driver.sv"
        `include "apb_reset_agent.sv"

        `include "apb_env.sv"
        `include "apb_test.sv"
    endpackage

/**********************************************************************************************************************
*  END OF FILE: apb_pkg.sv
*********************************************************************************************************************/